THERMO ALL
   200.000  1000.000  5000.000
! NASA Polynomial format for CHEMKIN-II
! see README file for disclaimer
AR                      AR  1               G    200.00   5000.00 1000.00      1
 2.50000000e+00 2.80607321e-14-2.32701659e-17 7.79829447e-21-9.11155357e-25    2
-7.45375000e+02 4.36600000e+00 2.50000000e+00-5.82136958e-14 1.06141476e-16    3
-7.84761333e-20 2.06574516e-23-7.45375000e+02 4.36600000e+00                   4
C                       C   1               G    200.00   5000.00 1000.00      1
 2.47498226e+00 8.64011929e-05-1.01325178e-07 4.64692686e-11-5.87731503e-15    2
 8.54573472e+04 4.89694985e+00 2.53378657e+00-1.48816040e-04 2.51500671e-07    3
-1.88747964e-10 5.29269932e-14 8.54455864e+04 4.61325305e+00                   4
C2H                     C   2H   1          G    200.00   5000.00 1000.00      1
 4.72139559e+00 1.32359549e-03 7.65068372e-07-5.14940019e-10 7.36354245e-14    2
 6.66006521e+04-1.71856069e+00 4.01925748e+00 4.13214795e-03-3.44776031e-06    3
 2.29361244e-09-6.28502689e-13 6.67410797e+04 1.66884983e+00                   4
C2H2                    C   2H   2          G    200.00   5000.00 1000.00      1
 5.02223749e+00 3.96264596e-03-8.20829533e-07-2.85649929e-11 1.98015842e-14    2
 2.56562780e+04-5.89796695e+00 1.44581772e+00 1.82683250e-02-2.22793481e-05    3
 1.42771141e-08-3.55661818e-12 2.63715620e+04 1.13561911e+01                   4
C2H3                    C   2H   3          G    200.00   5000.00 1000.00      1
 2.15349018e+00 1.22451457e-02-6.14404539e-06 1.48093889e-09-1.38213265e-13    2
 3.49009541e+04 1.24255790e+01 1.75610588e+00 1.38346829e-02-8.52835116e-06    3
 3.07047607e-09-5.35597560e-13 3.49804310e+04 1.43427285e+01                   4
C2H4                    C   2H   4          G    200.00   5000.00 1000.00      1
 2.32923141e-01 1.86761020e-02-9.80342021e-06 2.45377306e-09-2.35926437e-13    2
 5.53526916e+03 1.99773582e+01 1.37999702e+00 1.40878065e-02-2.92097694e-06    3
-2.13452246e-09 9.11147442e-13 5.30585438e+03 1.44433898e+01                   4
C2H5                    C   2H   5          G    200.00   5000.00 1000.00      1
 3.75894283e-01 2.09224709e-02-1.06843266e-05 2.60916612e-09-2.45815943e-13    2
 1.33794237e+04 2.19324486e+01 2.16625502e+00 1.37610279e-02 5.78378268e-08    3
-4.55227683e-09 1.54454479e-12 1.30213515e+04 1.32949930e+01                   4
C2H6                    C   2H   6          G    200.00   5000.00 1000.00      1
-9.39162113e-01 2.61720089e-02-1.34616992e-05 3.30289375e-09-3.12097942e-13    2
-1.07611305e+04 2.59063121e+01 1.82501487e+00 1.51153010e-02 3.12336270e-06    3
-7.75381417e-09 2.45207904e-12-1.13139659e+04 1.25707560e+01                   4
C3H7                    C   3H   7          G    250.00   3500.00 1000.00      1
 2.35156051e+00 2.74246855e-02-1.36908154e-05 3.35514575e-09-3.23981589e-13    2
 1.01707250e+04 1.35145484e+01-1.04791995e+00 4.10226074e-02-3.40876982e-05    3
 1.69530676e-08-3.72346205e-12 1.08506211e+04 2.99150765e+01                   4
C3H8                    C   3H   8          G    200.00   5000.00 1000.00      1
 9.20641409e-01 3.29494854e-02-1.66765872e-05 4.12359122e-09-4.00190440e-13    2
-1.41561236e+04 1.79356758e+01-1.21455954e+00 4.14902891e-02-2.94877929e-05    3
 1.26643950e-08-2.53539139e-12-1.37290834e+04 2.82367861e+01                   4
CH                      C   1H   1          G    200.00   5000.00 1000.00      1
 3.37627957e+00-1.21143157e-04 9.69465996e-07-3.89305903e-10 4.63620315e-14    2
 7.08445469e+04 2.80476100e+00 3.71486557e+00-1.47548716e-03 3.00098200e-06    3
-1.74364990e-09 3.84948031e-13 7.07768297e+04 1.17127927e+00                   4
CH2                     C   1H   2          G    200.00   5000.00 1000.00      1
 3.53245066e+00 2.20114905e-03-3.05697461e-07-8.62054079e-11 1.97651396e-14    2
 4.60440155e+04 2.63292262e+00 3.74382392e+00 1.35565598e-03 9.62542150e-07    3
-9.31698481e-10 2.31138408e-13 4.60017408e+04 1.61316879e+00                   4
CH2(S)                  C   1H   2          G    200.00   5000.00 1000.00      1
 2.64044175e+00 3.89119009e-03-1.43477007e-06 2.37240973e-10-1.39136758e-14    2
 5.08087160e+04 6.75114549e+00 4.21614957e+00-2.41164119e-03 8.01947685e-06    3
-6.06559031e-09 1.56179415e-12 5.04935744e+04-8.50733902e-01                   4
CH2CHO                  O   1H   3C   2     G    200.00   5000.00 1000.00      1
 2.94798131e+00 1.45651920e-02-7.49356762e-06 1.87044540e-09-1.82323244e-13    2
 1.55028604e+03 1.13619853e+01 2.69288424e+00 1.55855803e-02-9.02415004e-06    3
 2.89083367e-09-4.37420313e-13 1.60130545e+03 1.25926812e+01                   4
CH2CO                   C   2H   2O   1     G    200.00   5000.00 1000.00      1
 4.33729143e+00 9.33699691e-03-4.39637931e-06 9.88949688e-10-8.63225110e-14    2
-7.48311917e+03 1.59417110e+00 2.14047449e+00 1.81242647e-02-1.75772810e-05    3
 9.77621746e-09-2.28313945e-12-7.04375578e+03 1.21925430e+01                   4
CH2O                    H   2C   1O   1     G    200.00   5000.00 1000.00      1
 4.69195464e-01 1.20871438e-02-6.63394412e-06 1.70673325e-09-1.66860646e-13    2
-1.35701758e+04 2.05823651e+01 3.67988739e+00-7.55623875e-04 1.26302074e-05    3
-1.11360344e-08 3.04383128e-12-1.42123142e+04 5.09263257e+00                   4
CH2OH                   C   1H   3O   1     G    200.00   5000.00 1000.00      1
 3.44119170e+00 9.21164027e-03-4.18745102e-06 9.26308475e-10-8.05213258e-14    2
-3.16012376e+03 7.15745906e+00 3.42922492e+00 9.25950737e-03-4.25925167e-06    3
 9.74175574e-10-9.24881006e-14-3.15773040e+03 7.21519183e+00                   4
CH3                     C   1H   3          G    200.00   5000.00 1000.00      1
 2.76046463e+00 6.20364970e-03-2.20855773e-06 3.52842941e-10-1.98327525e-14    2
 1.66147681e+04 5.92182069e+00 3.58664806e+00 2.89891599e-03 2.74854284e-06    3
-2.95189077e-09 8.06350675e-13 1.64495314e+04 1.93596323e+00                   4
CH3CHO                  C   2H   4O   1     G    200.00   5000.00 1000.00      1
 9.96590574e-01 2.12592263e-02-1.13650710e-05 2.90734875e-09-2.87083467e-13    2
-2.10807853e+04 2.03188071e+01 2.46079397e+00 1.54024127e-02-2.57985059e-06    3
-2.94946485e-09 1.17711993e-12-2.13736260e+04 1.32548721e+01                   4
CH3O                    C   1H   3O   1     G    200.00   5000.00 1000.00      1
 5.74443531e-01 1.47199069e-02-7.74016881e-06 1.96701038e-09-1.94180320e-13    2
 1.23604905e+03 2.02217775e+01 1.49675601e+00 1.10306569e-02-2.20629394e-06    3
-1.72223954e-09 7.28132159e-13 1.05158655e+03 1.57721529e+01                   4
CH3OH                   C   1H   4O   1     G    200.00   5000.00 1000.00      1
-1.47987100e-01 1.84629596e-02-9.73380748e-06 2.45407041e-09-2.37706398e-13    2
-2.47427725e+04 2.48754627e+01 3.34423632e+00 4.49406590e-03 1.12195330e-05    3
-1.15148233e-08 3.25451702e-12-2.54412172e+04 8.02750340e+00                   4
CH4                     C   1H   4          G    200.00   5000.00 1000.00      1
-7.06145866e-01 1.51864609e-02-7.13580711e-06 1.67375885e-09-1.52892015e-13    2
-9.21994761e+03 2.26007083e+01 3.89942811e+00-3.23583504e-03 2.04976368e-05    3
-1.67485371e-08 4.45268196e-12-1.01410624e+04 3.81476172e-01                   4
CN                      C   1N   1          G    200.00   5000.00 1000.00      1
 2.71825043e+00 2.22309212e-03-1.30891267e-06 4.25346765e-10-4.97150090e-14    2
 5.18967469e+04 8.35827823e+00 3.66424500e+00-1.56088614e-03 4.36705473e-06    3
-3.35863150e-09 8.96279558e-13 5.17075480e+04 3.79440128e+00                   4
CO                      C   1O   1          G    200.00   5000.00 1000.00      1
 2.71449428e+00 2.05672640e-03-9.89797792e-07 2.26040507e-10-1.98121703e-14    2
-1.41503973e+04 7.82594967e+00 3.75251424e+00-2.09535342e-03 5.23832194e-06    3
-3.92603932e-09 1.01820779e-12-1.43580013e+04 2.81810342e+00                   4
CO2                     C   1O   2          G    200.00   5000.00 1000.00      1
 3.36612576e+00 5.46190472e-03-2.99036351e-06 7.63033672e-10-7.35465714e-14    2
-4.85877004e+04 4.93263369e+00 2.22771753e+00 1.00155377e-02-9.82081292e-06    3
 5.31666661e-09-1.21195481e-12-4.83600188e+04 1.04247954e+01                   4
H                       H   1               G    200.00   5000.00 1000.00      1
 2.50000000e+00 1.39443526e-12-3.97898542e-15 1.91753662e-18-2.67863269e-22    2
 2.54736599e+04-4.46682856e-01 2.50000000e+00 7.88907057e-12-1.37209384e-14    3
 8.41217193e-18-1.89152210e-21 2.54736599e+04-4.46682848e-01                   4
H2                      H   2               G    200.00   5000.00 1000.00      1
 4.00912475e+00-1.53371940e-03 1.62806503e-06-5.35274170e-10 5.97521864e-14    2
-1.17506714e+03-6.81731757e+00 3.00416922e+00 2.48610276e-03-4.40166821e-06    3
 3.48454799e-09-9.45203353e-13-9.74076035e+02-1.96898801e+00                   4
H2CN                    H   2C   1N   1     G    200.00   5000.00 1000.00      1
 2.04115515e+00 9.82901697e-03-5.41413427e-06 1.43096045e-09-1.45699967e-13    2
 2.87619167e+04 1.26601702e+01 2.31757391e+00 8.72334192e-03-3.75562169e-06    3
 3.25285399e-10 1.30718796e-13 2.87066330e+04 1.13266095e+01                   4
H2O                     H   2O   1          G    200.00   5000.00 1000.00      1
 3.46818930e+00 1.25793349e-03 5.11816268e-07-3.04627893e-10 3.95366379e-14    2
-3.01569447e+04 2.61200111e+00 4.13256435e+00-1.39956671e-03 4.49806656e-06    3
-2.96212809e-09 7.03911687e-13-3.02898197e+04-5.93224456e-01                   4
H2O2                    H   2O   2          G    200.00   5000.00 1000.00      1
 3.54004447e+00 6.32719048e-03-3.00091969e-06 7.22498370e-10-6.84279096e-14    2
-1.76596577e+04 6.25691155e+00 3.37370597e+00 6.99254447e-03-3.99895067e-06    3
 1.38785236e-09-2.34766406e-13-1.76263900e+04 7.05939864e+00                   4
HCCO                    H   1C   2O   1     G    200.00   5000.00 1000.00      1
 5.08985181e+00 5.18506807e-03-2.38092871e-06 5.23200438e-10-4.49225707e-14    2
 1.95240656e+04-9.90029958e-01 2.54746630e+00 1.53546101e-02-1.76352417e-05    3
 1.06927425e-08-2.58730808e-12 2.00325427e+04 1.12755105e+01                   4
HCCOH                   C   2O   1H   2     G    200.00   5000.00 1000.00      1
 6.23527496e+00 5.97008792e-03-1.87128565e-06 2.15511774e-10-2.49832022e-15    2
 7.18589540e+03-9.20691740e+00 2.74316416e+00 1.99385311e-02-2.28239504e-05    3
 1.41839550e-08-3.49460912e-12 7.88431756e+03 7.64049858e+00                   4
HCN                     H   1C   1N   1     G    200.00   5000.00 1000.00      1
 3.74782550e+00 3.19046862e-03-1.05704758e-06 1.55362727e-10-7.85766702e-15    2
 1.44399459e+04 1.90733211e+00 2.48224378e+00 8.25279549e-03-8.65053789e-06    3
 5.21768960e-09-1.27343938e-12 1.46930622e+04 8.01303233e+00                   4
HCNN                    C   1N   2H   1     G    200.00   5000.00 1000.00      1
 4.98981658e+00 5.89302215e-03-2.99250038e-06 7.19510963e-10-6.67290488e-14    2
 5.37733729e+04-1.89753630e-01 2.53645525e+00 1.57064675e-02-1.77126684e-05    3
 1.05329563e-08-2.52009038e-12 5.42640451e+04 1.16462966e+01                   4
HCNO                    H   1N   1C   1O   1G    200.00   5000.00 1000.00      1
 4.04560456e+00 7.87589814e-03-4.37486726e-06 1.12800925e-09-1.10378868e-13    2
 1.89953177e+04 3.83002454e+00 2.38041291e+00 1.45366647e-02-1.43660172e-05    3
 7.78877585e-09-1.77557052e-12 1.93283560e+04 1.18636117e+01                   4
HCO                     H   1C   1O   1     G    200.00   5000.00 1000.00      1
 2.16910758e+00 6.28662528e-03-3.49267468e-06 9.06066457e-10-8.86584634e-14    2
 4.21405817e+03 1.30418141e+01 3.89571999e+00-6.19824377e-04 6.86699980e-06    3
-6.00038320e-09 1.63795395e-12 3.86873569e+03 4.71190730e+00                   4
HNCO                    H   1N   1C   1O   1G    200.00   5000.00 1000.00      1
 3.41508897e+00 8.63397044e-03-4.86846097e-06 1.27978182e-09-1.27386717e-13    2
-1.55617480e+04 7.12400489e+00 3.42344553e+00 8.60054423e-03-4.81832165e-06    3
 1.24635560e-09-1.19030164e-13-1.55634193e+04 7.08368935e+00                   4
HNO                     H   1N   1O   1     G    200.00   5000.00 1000.00      1
 2.47117866e+00 4.71558439e-03-1.76366752e-06 3.76611743e-10-3.67093701e-14    2
 1.19016409e+04 1.12866703e+01 3.99629668e+00-1.38488771e-03 7.38704062e-06    3
-5.72386035e-09 1.48840865e-12 1.15966173e+04 3.92885746e+00                   4
HO2                     H   1O   2          G    200.00   5000.00 1000.00      1
 3.02157955e+00 4.45643776e-03-2.32743819e-06 6.49879149e-10-7.07552917e-14    2
 4.41857297e+02 9.12939911e+00 3.34788125e+00 3.15123095e-03-3.69627964e-07    3
-6.55327666e-10 2.55546412e-13 3.76596957e+02 7.55518201e+00                   4
HOCN                    H   1N   1C   1O   1G    200.00   5000.00 1000.00      1
 3.72572353e+00 7.23598680e-03-3.85095113e-06 9.61231844e-10-9.18441695e-14    2
-2.81954060e+03 5.89630053e+00 3.73205550e+00 7.21065888e-03-3.81295926e-06    3
 9.35903928e-10-8.55121907e-14-2.82080699e+03 5.86575239e+00                   4
N                       N   1               G    200.00   5000.00 1000.00      1
 2.49388718e+00 1.03463806e-05 1.86374207e-09-6.88831219e-12 2.02531990e-15    2
 5.61062724e+04 4.22664607e+00 2.50529382e+00-3.52801781e-05 7.03035801e-08    3
-5.25148709e-11 1.34319596e-14 5.61039911e+04 4.17161563e+00                   4
N2                      N   2               G    200.00   5000.00 1000.00      1
 2.83503116e+00 1.62289122e-03-6.35527663e-07 1.14074754e-10-7.55177506e-15    2
-8.79411301e+02 6.50778052e+00 3.77288186e+00-2.12851156e-03 4.99157651e-06    3
-3.63732803e-09 9.30298921e-13-1.06698144e+03 1.98319304e+00                   4
N2O                     N   2O   1          G    200.00   5000.00 1000.00      1
 3.73479390e+00 4.92113121e-03-2.64141316e-06 6.75980188e-10-6.61702123e-14    2
 8.45788432e+03 3.70529797e+00 2.32814401e+00 1.05477307e-02-1.10813125e-05    3
 6.30257972e-09-1.47282010e-12 8.73921430e+03 1.04915705e+01                   4
NCO                     N   1C   1O   1     G    200.00   5000.00 1000.00      1
 3.74927426e+00 5.30790964e-03-3.10805898e-06 8.36757922e-10-8.48886664e-14    2
 1.44911854e+04 5.04715208e+00 2.72689023e+00 9.39744577e-03-9.24236316e-06    3
 4.92629404e-09-1.10727270e-12 1.46956622e+04 9.97956404e+00                   4
NH                      N   1H   1          G    200.00   5000.00 1000.00      1
 3.35038855e+00 7.69069409e-05 5.26492144e-07-2.20841683e-10 2.78388685e-14    2
 4.19316590e+04 2.69488024e+00 3.70656804e+00-1.34781103e-03 2.66356910e-06    3
-1.64555966e-09 3.84018362e-13 4.18604231e+04 9.76520072e-01                   4
NH2                     N   1H   2          G    200.00   5000.00 1000.00      1
 2.95847561e+00 2.91131160e-03-6.98110918e-07 6.04794113e-11 8.01681473e-16    2
 2.21350150e+04 5.86712912e+00 4.21525850e+00-2.11581995e-03 6.84258639e-06    3
-4.96665213e-09 1.25758457e-12 2.18836585e+04-1.96121809e-01                   4
NH3                     N   1H   3          G    200.00   5000.00 1000.00      1
 2.21298890e+00 6.60936780e-03-2.45237546e-06 4.68872021e-10-3.84533357e-14    2
-6.40566075e+03 8.82653479e+00 3.61275208e+00 1.01031508e-03 5.94620362e-06    3
-5.13018070e-09 1.36130984e-12-6.68561338e+03 2.07348658e+00                   4
NNH                     N   2H   1          G    200.00   5000.00 1000.00      1
 2.54113032e+00 5.56550055e-03-3.05549572e-06 7.98506858e-10-8.00621699e-14    2
 2.90670769e+04 1.10772085e+01 3.58561560e+00 1.38755945e-03 3.21141594e-06    3
-3.37943425e-09 9.64423106e-13 2.88581799e+04 6.03817085e+00                   4
NO                      N   1O   1          G    200.00   5000.00 1000.00      1
 2.59342250e+00 2.64431541e-03-1.52126173e-06 4.10437136e-10-4.18290559e-14    2
 1.01478971e+04 9.96666481e+00 4.01175979e+00-3.02903373e-03 6.98876198e-06    3
-5.26291200e-09 1.37650823e-12 9.86422962e+03 3.12400729e+00                   4
NO2                     N   1O   2          G    200.00   5000.00 1000.00      1
 2.81928779e+00 6.66768263e-03-4.20601268e-06 1.21236074e-09-1.27472090e-13    2
 3.01997274e+03 1.10216145e+01 3.02085922e+00 5.86139688e-03-2.99658406e-06    3
 4.06074994e-10 7.40993455e-14 2.97965845e+03 1.00491489e+01                   4
O                       O   1               G    200.00   5000.00 1000.00      1
 2.51192991e+00 5.18142381e-05-6.87799798e-08 2.62748075e-11-2.94338252e-15    2
 2.92348465e+04 5.08799277e+00 3.00827493e+00-1.93356585e-03 2.90929014e-06    3
-1.95910528e-09 4.93401638e-13 2.91355775e+04 2.69341496e+00                   4
O2                      O   2               G    200.00   5000.00 1000.00      1
 2.60925233e+00 2.97662855e-03-1.89478508e-06 5.67712477e-10-6.16566842e-14    2
-8.64566737e+02 9.06957329e+00 3.45703182e+00-4.14489410e-04 3.19189186e-06    3
-2.82340548e-09 7.86122806e-13-1.03412263e+03 4.97952732e+00                   4
OH                      O   1H   1          G    200.00   5000.00 1000.00      1
 3.57809111e+00-5.01489805e-04 9.11030475e-07-3.31737105e-10 3.86587420e-14    2
 3.69246914e+03 1.85722061e+00 3.96510000e+00-2.04952537e-03 3.23308382e-06    3
-1.87977267e-09 4.25667633e-13 3.61506736e+03-9.87357253e-03                   4
END
